

  



  







             






 
  
  
   
 








 






 






 







 



 


 





 


          







 



 


 





 


          




























         




 




 




  












             











































































































               









  


























********















****************





    















































***********************************************************************************

 

 

 

 













































































































    
   










        









    
   










        ******   **********



























************************

















*****************************************************************************************************************************************************************************************************


																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			   																																																																																																																																																																																																																																																																																																																																		             																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								 																																																																																																																																																																																																																																																																																																																																																																																																																																											 																																						     																																												            																																																												    																																																																																																																																																																																																																			    																																																																																																																																								  															   		   																							   																																																		      									     																				         																																																																																																																																																																																																																																																																																								        																																																										       																																																																																																																																																																																																																																											   																									   			 																																																																																																																																																																																																										   																																																																																																																																																																																																																																																																														                         																																																																																																																																																																																																																																																																																																																											        																																																																																																																																																																																																																																																																																																																																																																																																																	   																																																																																																																																																																																																																																																																																																																							    																																																																																																																																																																																																																																																																																																																																																																																																													                              																																		  																														   						                                                                                                                                                                                                                																								  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																									 																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																						                                                                                                                                                                                                                                                                                                                              .....................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                             .....................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  